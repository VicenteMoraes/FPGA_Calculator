library verilog;
use verilog.vl_types.all;
entity pre_projeto_vlg_vec_tst is
end pre_projeto_vlg_vec_tst;
