library verilog;
use verilog.vl_types.all;
entity bcd_converter_vlg_vec_tst is
end bcd_converter_vlg_vec_tst;
